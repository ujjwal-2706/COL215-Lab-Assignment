----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/14/2022 02:57:25 PM
-- Design Name: 
-- Module Name: comparator - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity comparator is
  Port ( 
    comparator_enable : in std_logic;
    input1 : inout signed(15 downto 0) := x"ffff";
    input2 : in signed(15 downto 0);
    address : inout integer := 0;
    index : in integer
  );
end comparator;

architecture Behavioral of comparator is

begin
input1 <= input2 when ((input1 < input2) and (comparator_enable = '1')) else input1;
address <= index when ((input1 < input2) and (comparator_enable = '1')) else address;
end Behavioral;
